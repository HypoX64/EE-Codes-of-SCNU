LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY timectr_clkdiv IS
	PORT(
		sysclk:IN STD_LOGIC;
		clk_01:OUT STD_LOGIC);
	END ENTITY timectr_clkdiv;
	
ARCHITECTURE rt1 OF timectr_clkdiv IS
SIGNAL div1:STD_LOGIC_VECTOR(3 DOWNTO 0):="0000";--divide by 256counter
SIGNAL div2:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000"; --10
SIGNAL div3:STD_LOGIC_VECTOR(7 DOWNTO 0):="00"; --3
SIGNAL clk1,clk2:STD_LOGIC;

BEGIN
div_10:PROCESS(clk1)IS
BEGIN